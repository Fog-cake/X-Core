// Copyright 2015 ETH Zurich and University of Bologna.
// Copyright 2017 Embecosm Limited <www.embecosm.com>
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.

/*module dp_ram
  #(
    parameter ADDR_WIDTH = 34
  )(
    // Clock and Reset
    input  logic clk,

    input  logic                   en_a_i,
    input  logic [ADDR_WIDTH-1:0]  addr_a_i,
    input  logic [31:0]            wdata_a_i,
    output logic [127:0]           rdata_a_o,
    input  logic                   we_a_i,
    input  logic [3:0]             be_a_i,

    input  logic                   en_b_i,
    input  logic [ADDR_WIDTH-1:0]  addr_b_i,
    input  logic [31:0]            wdata_b_i,
    output logic [31:0]            rdata_b_o,
    input  logic                   we_b_i,
    input  logic [3:0]             be_b_i,
	output logic 					cmd_ready
  );



  localparam bytes = 2**20;//ADDR_WIDTH;

  reg   [7:0] mem[0:bytes-1];
  logic [19:0] addr_b_int;

  initial begin
    $readmemh("F:/riscv_dbg_201808010/dhrystone.verilog", mem); 
  end

  always_comb addr_b_int = {addr_b_i[31:2], 2'b0};

  always @(posedge clk)
  begin

    rdata_a_o[  0+: 8] <= mem[addr_a_i +  0];
    rdata_a_o[  8+: 8] <= mem[addr_a_i +  1];
    rdata_a_o[ 16+: 8] <= mem[addr_a_i +  2];
    rdata_a_o[ 24+: 8] <= mem[addr_a_i +  3];
    rdata_a_o[ 32+: 8] <= mem[addr_a_i +  4];
    rdata_a_o[ 40+: 8] <= mem[addr_a_i +  5];
    rdata_a_o[ 48+: 8] <= mem[addr_a_i +  6];
    rdata_a_o[ 56+: 8] <= mem[addr_a_i +  7];
    rdata_a_o[ 64+: 8] <= mem[addr_a_i +  8];
    rdata_a_o[ 72+: 8] <= mem[addr_a_i +  9];
    rdata_a_o[ 80+: 8] <= mem[addr_a_i + 10];
    rdata_a_o[ 88+: 8] <= mem[addr_a_i + 11];
    rdata_a_o[ 96+: 8] <= mem[addr_a_i + 12];
    rdata_a_o[104+: 8] <= mem[addr_a_i + 13];
    rdata_a_o[112+: 8] <= mem[addr_a_i + 14];
    rdata_a_o[120+: 8] <= mem[addr_a_i + 15];

    //* addr_b_i is the actual memory address referenced 
cmd_ready <= 0;
    if (en_b_i)
    begin
      //* handle writes 
	  cmd_ready <= 1;
      if (we_b_i)
      begin
        if (be_b_i[0]) mem[addr_b_int    ] <= wdata_b_i[ 0+:8];
        if (be_b_i[1]) mem[addr_b_int + 1] <= wdata_b_i[ 8+:8];
        if (be_b_i[2]) mem[addr_b_int + 2] <= wdata_b_i[16+:8];
        if (be_b_i[3]) mem[addr_b_int + 3] <= wdata_b_i[24+:8];
      end
      //* handle reads 
      else
      begin
        rdata_b_o[ 7: 0] <= mem[addr_b_int    ];
        rdata_b_o[15: 8] <= mem[addr_b_int + 1];
        rdata_b_o[23:16] <= mem[addr_b_int + 2];
        rdata_b_o[31:24] <= mem[addr_b_int + 3];
      end
    end
	else
		cmd_ready <= 0;
  end

  function [7:0] readByte;
    //verilator public 
    input integer byte_addr;
    readByte = mem[byte_addr];
  endfunction

  task writeByte;
    // verilator public 
    input integer byte_addr;
    input [7:0] val;
    mem[byte_addr] = val;
  endtask

endmodule*/
// Copyright 2015 ETH Zurich and University of Bologna.
// Copyright 2017 Embecosm Limited <www.embecosm.com>
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.

module dp_ram
  #(
    parameter ADDR_WIDTH = 34
  )(
    // Clock and Reset
    input  logic 					clk,
	input  logic					rst_n,
    input  logic                   	en_a_i,
    input  logic [ADDR_WIDTH-1:0]  	addr_a_i,
    input  logic [31:0]            	wdata_a_i,
    output logic [127:0]          	rdata_a_o,
    input  logic                   	we_a_i,
    input  logic [3:0]             	be_a_i,

    input  logic                   	en_b_i,
    input  logic [ADDR_WIDTH-1:0]  	addr_b_i,
    input  logic [31:0]            	wdata_b_i,
    output logic [31:0]            	rdata_b_o,
    input  logic                   	we_b_i,
    input  logic [3:0]             	be_b_i,
	output logic 					cmd_ready
  );



  localparam bytes = 2**20;//ADDR_WIDTH;

  reg   [7:0] mem[0:bytes-1];
  logic [19:0] addr_b_int;

   //initial begin
   // $readmemh("C:/Users/PerfxLab-ChenBotao/Desktop/e200_opensource-master/riscv-tools/riscv-tests/isa/generated/rv32ui-p-add.verilog", mem); 
   //end

  always_comb addr_b_int = {addr_b_i[31:2], 2'b0};

  always @(posedge clk )
//	if (!rst_n)
//		begin
//			mem[0] <= 8'H97;
//			mem[1] <= 8'H22;
//			mem[2] <= 8'H01;
//			mem[3] <= 8'He0;
//			mem[4] <= 8'H13;
//			mem[5] <= 8'H02;
//			mem[6] <= 8'Hc0;
//			mem[7] <= 8'H9e;
//			mem[8] <= 8'H33;
//			mem[9] <= 8'H03;
//			mem[10] <= 8'H52;
//			mem[11] <= 8'H00;
//			mem[12] <= 8'H93;
//			mem[13] <= 8'H03;
//			mem[14] <= 8'Hf0;
//			mem[15] <= 8'H06;
//			mem[16] <= 8'H23;
//			mem[17] <= 8'H20;
//			mem[18] <= 8'H73;
//			mem[19] <= 8'H00;
//			mem[20] <= 8'H67;
//			mem[21] <= 8'H80;
//			mem[22] <= 8'Hc2;
//			mem[23] <= 8'H9e;
//			mem[24] <= 8'H6f;
//			mem[25] <= 8'H00;
//			mem[26] <= 8'H00;
//			mem[27] <= 8'H00;
//			mem[28] <= 8'H6f;
//			mem[29] <= 8'H00;
//			mem[30] <= 8'H00;
//			mem[31] <= 8'H00;	
			
//		end
//	else
	  begin

		rdata_a_o[  0+: 8] <= mem[addr_a_i +  0];
		rdata_a_o[  8+: 8] <= mem[addr_a_i +  1];
		rdata_a_o[ 16+: 8] <= mem[addr_a_i +  2];
		rdata_a_o[ 24+: 8] <= mem[addr_a_i +  3];
		rdata_a_o[ 32+: 8] <= mem[addr_a_i +  4];
		rdata_a_o[ 40+: 8] <= mem[addr_a_i +  5];
		rdata_a_o[ 48+: 8] <= mem[addr_a_i +  6];
		rdata_a_o[ 56+: 8] <= mem[addr_a_i +  7];
		rdata_a_o[ 64+: 8] <= mem[addr_a_i +  8];
		rdata_a_o[ 72+: 8] <= mem[addr_a_i +  9];
		rdata_a_o[ 80+: 8] <= mem[addr_a_i + 10];
		rdata_a_o[ 88+: 8] <= mem[addr_a_i + 11];
		rdata_a_o[ 96+: 8] <= mem[addr_a_i + 12];
		rdata_a_o[104+: 8] <= mem[addr_a_i + 13];
		rdata_a_o[112+: 8] <= mem[addr_a_i + 14];
		rdata_a_o[120+: 8] <= mem[addr_a_i + 15];

		/* addr_b_i is the actual memory address referenced */
		cmd_ready <= 0;
		if (en_b_i)
		begin
		  /* handle writes */
		  cmd_ready <= 1;
		  if (we_b_i)
		  begin
			if (be_b_i[0]) mem[addr_b_int    ] <= wdata_b_i[ 0+:8];
			if (be_b_i[1]) mem[addr_b_int + 1] <= wdata_b_i[ 8+:8];
			if (be_b_i[2]) mem[addr_b_int + 2] <= wdata_b_i[16+:8];
			if (be_b_i[3]) mem[addr_b_int + 3] <= wdata_b_i[24+:8];
		  end
		  /* handle reads */
		  else
		  begin
			rdata_b_o[ 7: 0] <= mem[addr_b_int    ];
			rdata_b_o[15: 8] <= mem[addr_b_int + 1];
			rdata_b_o[23:16] <= mem[addr_b_int + 2];
			rdata_b_o[31:24] <= mem[addr_b_int + 3];
		  end
		end
		else
			cmd_ready <= 0;
	  end

	  function [7:0] readByte;
		/* verilator public */
		input integer byte_addr;
		readByte = mem[byte_addr];
	  endfunction

  task writeByte;
    /* verilator public */
    input integer byte_addr;
    input [7:0] val;
    mem[byte_addr] = val;
  endtask

endmodule



